//***********************************************************************
//    Copyright (c) 2024 @freecity
//    All Rights Reserved.
//***********************************************************************
//-----------------------------------------------------------------------
// File:        cbb_ecc_enc.v
// Auther:      churchmice ( firefoxelectric@gmail.com )
// Created:     17:07:04, May 19, 2024
//-----------------------------------------------------------------------
// Abstract:    Haming code + extra parity that could correct one bit error
//              and detect 2 bits error. Maximal user data length is 256 bits
//              The error injection function is used to test the system behavior
//              when an ecc error occurs
//parity bits   data bits   total bits
//2             1           3
//3             4           7
//4             11          15
//5             26          31
//6             57          63
//7             120         127
//8             247         255
//9             502         511
`ifndef __CBB_ECC_ENC__
`define __CBB_ECC_ENC__
module cbb_ecc_enc #(
    parameter   DW = 32,
    parameter   EW = 7      //shall set accordingly to the DW length, shall include an extra bit for the overall parity
)(
    input   wire                clk,
    input   wire                rst_n,
    input   wire                inj_1bit_err,   //to inject single bit error
    input   wire                inj_2bit_err,   //to inject double bit error
    input   wire [DW-1:0]       din,
    output  reg  [DW+EW-1:0]    dout
);
    //define the maximal generation matrix
    wire [255:0] g_matrix [8:0];
    wire [EW-1:0] ecc;
    assign  g_matrix[00] = 256'b1010101011010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101101010101010101010101010101010101010101010101010101010101010101101010101010101010101010101010110101010101010110101011011;
    assign  g_matrix[01] = 256'b0011001101100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110110011001100110011001100110011001100110011001100110011001100110110011001100110011001100110011011001100110011011001101101;
    assign  g_matrix[02] = 256'b0011110001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000111100001111000011110000111100001111000011110000111100001111000111100001111000011110000111100011110000111100011110001110;
    assign  g_matrix[03] = 256'b1100000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000111111110000000011111111000000001111111100000000111111110000000111111110000000011111111000000011111111000000011111110000;
    assign  g_matrix[04] = 256'b0000000001111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111000000000000000111111111111111100000000000000001111111111111111000000000000000111111111111111100000000000000011111111111111100000000000;
    assign  g_matrix[05] = 256'b0000000001111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000111111111111111111111111111111100000000000000000000000000;
    assign  g_matrix[06] = 256'b0000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000;
    assign  g_matrix[07] = 256'b0000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign  g_matrix[08] = 256'b1111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

    generate 
        for ( genvar g = 0 ; g < EW - 1 ; g ++ ) begin: gen_ecc
            assign ecc[g] = ^(din & g_matrix[g][DW-1:0]) ;
        end
    endgenerate

    //extra bit for the SECDED
    assign  ecc[EW-1] = ^{ ecc[0+:EW-1], din};

    always @(posedge clk or negedge rst_n ) begin
        if ( ~rst_n ) begin
            dout    <= {(DW+EW){1'b0}};
        end
        //note, we only need to generate an error
        else if ( inj_1bit_err ) begin
            dout    <= { ecc, din[DW-1:1], ~din[0] };
        end
        else if ( inj_2bit_err ) begin
            dout    <= { ecc[EW-1:1],~ecc[0], din[DW-1:1], ~din[0] };
        end
        else begin
            dout    <= { ecc, din };
        end
    end
endmodule
`endif
//-----------------------------------------------------------------------
// Local Variables:
// verilog-library-directories:()
// End:

